library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity InstructionMemory is
	port (
		ADDRESS: in STD_LOGIC_VECTOR (31 downto 0);
		DATA: out STD_LOGIC_VECTOR (31 downto 0)
	);
end InstructionMemory;


architecture Behavioral of InstructionMemory is	  

    type MemoryArray is array(0 to 63) of STD_LOGIC_VECTOR (31 downto 0);
    signal instrMemory: MemoryArray := (
        "00000000000000000100000000100101",
        "10001100000011010000000000110000",
        "10001100000110000000000000110100",
        "10001100000110010000000000111000",
        "00000000000110000101000000100000",
        "10101101000010100000000000000000",
        "10101101000010100000000000000100",
        "00000001101110000100100000100010",
        "00000001001110000100100000100010",
        "10001101000010110000000000000000",
         "10001101000011000000000000000100",
         "00000001011011000101000000100000",
         "10101101000010100000000000001000",
         "00000001000110010100000000100000",
         "00000001001110000100100000100010",
         "00000000000010010000100000101010",
         "00010000001000000000000000000001",
         "00001000000000000000000000001001",
         "00000000000001000010000000100100",
         "00000000000011010010100000100000",
         "00001000000000000000000000010110",
         "00000000000110001000000000100010",
         "00000001000000000100000000100100",
         "00000001000010000100100000100000",
         "00000001001010010100100000100000",
         "00000000100010010101000000100000",
         "10001101010100000000000000000000",
         "00000001000110000100000000100000",
         "00000001000001010000100000101010",
         "00010100001000001111111111111001",
         "00000000000000001100000000100111",
         "00000010000110001000000000100111",
         "00001000000000000000000000010101",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX",
         "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX"
    );

    begin
	 
    DATA <= instrMemory(to_integer(unsigned(ADDRESS)) / 4 );

end Behavioral;